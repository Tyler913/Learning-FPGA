module TouchButton_LED(
    input wire system_clock,
    input wire system_reset_n,
    input wire touch_button,

    output reg led
);

reg touch_key_1;
reg touch_key_2;
reg touch_flag;



endmodule
